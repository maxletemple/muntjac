`ifndef MUNTJAC_METADATA_TABLE_UTIL_SVH
`define MUNTJAC_METADATA_TABLE_UTIL_SVH

`define MUNTJAC_TRANSITION_TABLE_INIT_STATE 8'h00

`endif 